
module add_lower_bytes(    
    input a[3:0], b[3:0]
    output c, v[3:0]

);

endmodule;



module toplevel(
    input a[7:0], b[7:0], sub    
    output o[7:0]


);



endmodule;
